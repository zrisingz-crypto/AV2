//==============================================================================
// Real Coefficient Decoder Module for AV2
// Implements token parsing, run-length decoding, and EOB processing
//==============================================================================

`timescale 1ns / 1ps

// Note: This module uses internal memory for coefficients to comply with Verilog standards
// External modules should handle the unpacked array interface differently
module av2_coeff_decoder_real #(
    parameter MAX_COEFFS = 4096,
    parameter MAX_TX_SIZE = 64
)(
    input  wire                      clk,
    input  wire                      rst_n,
    
    // Input from entropy decoder
    input  wire [15:0]              context_idx,
    input  wire [15:0]              context_prob,
    input  wire [15:0]              decoded_symbol,
    input  wire                      symbol_valid,
    output reg                       symbol_ready,
    
    // Output coefficients - individual access
    output reg  signed [15:0]       coeff_out,
    output reg  [11:0]              coeff_addr,
    output reg                       coeff_valid,
    input  wire                      coeff_ready,
    
    // Output control
    output reg  [15:0]              num_coeffs,
    output reg                       coeffs_valid,
    input  wire                      coeffs_ready,
    
    // Transform parameters
    input  wire [5:0]               tx_size,
    input  wire [3:0]               tx_type,
    input  wire [7:0]               qindex,
    
    // Control
    input  wire                      start,
    output wire                      done
);

// Internal memory for coefficients
reg signed [15:0] coeffs [0:MAX_COEFFS-1];

// State machine
localparam IDLE       = 3'd0;
localparam TOKEN_PARSE = 3'd1;
localparam COEFF_GEN   = 3'd2;
localparam RUN_LENGTH = 3'd3;
localparam EOB_CHECK   = 3'd4;
localparam OUTPUT     = 3'd5;
localparam DONE       = 3'd6;

reg [2:0] state, state_next;

// Processing registers
reg [15:0] symbol_buf;
reg        symbol_buf_valid;
reg [11:0] coeff_idx;
reg [11:0] zero_run_count;
reg [11:0] processed_coeffs;
reg [15:0] eob_pos;
reg        eob_found;
reg [4:0]  scan_pos;
reg [15:0] last_nonzero_pos;

// Constants for scan orders
// Simplified 4x4 scan order (zigzag-like)
wire [4:0] scan_order_4x4 [0:15];
assign scan_order_4x4[0] = 5'd0;   // [0,0]
assign scan_order_4x4[1] = 5'd1;   // [1,0]
assign scan_order_4x4[2] = 5'd4;   // [0,1]
assign scan_order_4x4[3] = 5'd8;   // [0,2]
assign scan_order_4x4[4] = 5'd5;   // [1,1]
assign scan_order_4x4[5] = 5'd2;   // [2,0]
assign scan_order_4x4[6] = 5'd3;   // [3,0]
assign scan_order_4x4[7] = 5'd6;   // [2,1]
assign scan_order_4x4[8] = 5'd9;   // [1,2]
assign scan_order_4x4[9] = 5'd12;  // [1,3]
assign scan_order_4x4[10] = 5'd13; // [0,3]
assign scan_order_4x4[11] = 5'd14; // [0,4]
assign scan_order_4x4[12] = 5'd10; // [2,2]
assign scan_order_4x4[13] = 5'd7;  // [3,1]
assign scan_order_4x4[14] = 5'd11; // [3,2]
assign scan_order_4x4[15] = 5'd15; // [2,3]

// For larger transforms, we'll use a simplified row-major scan
reg [4:0] current_scan_pos;
reg [11:0] max_coeffs;

integer i;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
        symbol_ready <= 1'b0;
        coeffs_valid <= 1'b0;
        coeff_idx <= 12'd0;
        zero_run_count <= 12'd0;
        processed_coeffs <= 12'd0;
        eob_pos <= 16'd0;
        eob_found <= 1'b0;
        symbol_buf <= 16'd0;
        symbol_buf_valid <= 1'b0;
        last_nonzero_pos <= 16'd0;
        current_scan_pos <= 5'd0;
        coeff_out <= 16'sd0;
        coeff_addr <= 12'd0;
        coeff_valid <= 1'b0;
        
        for (i = 0; i < MAX_COEFFS; i = i + 1) begin
            coeffs[i] <= 16'sd0;
        end
        
        num_coeffs <= 16'd0;
    end else begin
        state <= state_next;
        
        case (state)
            IDLE: begin
                coeffs_valid <= 1'b0;
                coeff_valid <= 1'b0;
                symbol_ready <= 1'b0;
                eob_found <= 1'b0;
                coeff_idx <= 12'd0;
                processed_coeffs <= 12'd0;
                zero_run_count <= 12'd0;
                last_nonzero_pos <= 16'd0;
                
                if (start) begin
                    // Determine max coefficients based on transform size
                    case (tx_size)
                        6'd4:  max_coeffs <= 12'd16;
                        6'd8:  max_coeffs <= 12'd64;
                        6'd16: max_coeffs <= 12'd256;
                        6'd32: max_coeffs <= 12'd1024;
                        6'd64: max_coeffs <= 12'd4096;
                        default: max_coeffs <= 12'd256;  // Default to 16x16
                    endcase
                    
                    state <= TOKEN_PARSE;
                    symbol_ready <= 1'b1;
                end
            end
            
            TOKEN_PARSE: begin
                // Read symbols from entropy decoder and parse coefficients
                if (symbol_valid && symbol_ready) begin
                    $display("[TIME %0t] Coefficient decoder: received symbol %d from entropy decoder", $time, decoded_symbol);
                    
                    // Parse symbol to coefficient
                    // Simplified parsing: symbol value directly becomes coefficient
                    // In full implementation, this would use token tables
                    
                    // Check for EOB (End of Block) - symbol 65535 indicates EOB
                    if (decoded_symbol == 16'hFFFF) begin
                        eob_found <= 1'b1;
                        $display("[TIME %0t] Coefficient decoder: EOB found at position %d", $time, coeff_idx);
                        state <= OUTPUT;
                    end else if (coeff_idx < max_coeffs) begin
                        // Store coefficient
                        coeffs[coeff_idx] <= decoded_symbol;
                        
                        // Track last non-zero position
                        if (decoded_symbol != 16'sd0) begin
                            last_nonzero_pos <= coeff_idx;
                        end
                        
                        coeff_idx <= coeff_idx + 1;
                        
                        // Request next symbol
                        symbol_ready <= 1'b1;
                        
                        // Check if we've reached max coefficients
                        if (coeff_idx >= max_coeffs - 1) begin
                            state <= OUTPUT;
                        end
                    end else begin
                        // Reached max coefficients without EOB
                        state <= OUTPUT;
                    end
                end else if (!symbol_valid) begin
                    // Wait for entropy decoder to provide symbol
                    symbol_ready <= 1'b1;
                end
            end
            
            // These states are not needed in the simplified implementation
            // They can be added later for full token parsing support
            
            EOB_CHECK: begin
                // Check for End of Block
                // Simplified: if we've processed enough coefficients or received EOB signal
                if (coeff_idx >= max_coeffs || eob_found) begin
                    eob_pos <= last_nonzero_pos;
                    state <= OUTPUT;
                end else begin
                    state <= TOKEN_PARSE;  // Continue parsing
                    symbol_ready <= 1'b1;
                end
            end
            
            OUTPUT: begin
                // Prepare output
                coeffs_valid <= 1'b1;
                num_coeffs <= last_nonzero_pos + 1;  // Number of coefficients up to last non-zero
                
                // Output coefficients one by one
                if (coeffs_valid && !coeff_valid) begin
                    coeff_addr <= 12'd0;
                    coeff_out <= coeffs[0];
                    coeff_valid <= 1'b1;
                    $display("[TIME %0t] Coefficient decoder: Starting output, num_coeffs=%0d, last_nonzero=%0d", 
                             $time, num_coeffs, last_nonzero_pos);
                end else if (coeff_valid && coeff_ready && coeff_addr < num_coeffs-1) begin
                    coeff_addr <= coeff_addr + 1;
                    coeff_out <= coeffs[coeff_addr + 1];
                end else if (coeff_valid && coeff_ready && coeff_addr >= num_coeffs-1) begin
                    coeff_valid <= 1'b0;
                    coeffs_valid <= 1'b0;
                    $display("[TIME %0t] Coefficient decoder: All %0d coefficients output, moving to DONE", 
                             $time, num_coeffs);
                    state <= DONE;
                end
                
                // Also allow external ready signal to trigger completion
                if (coeffs_ready) begin
                    coeffs_valid <= 1'b0;
                    state <= DONE;
                end
            end
            
        DONE: begin
            coeffs_valid <= 1'b0;
            coeff_valid <= 1'b0;
            symbol_ready <= 1'b0;
            state <= IDLE;
        end
            
            default: begin
                state <= IDLE;
            end
        endcase
    end
end

// State transition logic
always @(*) begin
    state_next = state;
    
    case (state)
        IDLE: begin
            if (start)
                state_next = TOKEN_PARSE;
        end
        
        TOKEN_PARSE: begin
            // Stay in TOKEN_PARSE until EOB found or max coeffs reached
            if (eob_found || coeff_idx >= max_coeffs)
                state_next = OUTPUT;
        end
        
        OUTPUT: begin
            // Automatically transition to DONE after outputting all coefficients
            // Don't wait for coeffs_ready - it's optional
            if (coeff_valid && coeff_ready && coeff_addr >= num_coeffs-1)
                state_next = DONE;
            else if (coeffs_ready)
                state_next = DONE;
        end
        
        DONE: begin
            state_next = IDLE;
        end
        
        default: begin
            state_next = IDLE;
        end
    endcase
end

assign done = (state == DONE);

endmodule
